--
-- Copyright (C) 2021 Kiran Dsouza. All rights reserved.
-- 

